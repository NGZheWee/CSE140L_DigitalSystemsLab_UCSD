library verilog;
use verilog.vl_types.all;
entity display_tb_file_sv_unit is
end display_tb_file_sv_unit;
