library verilog;
use verilog.vl_types.all;
entity design_sv_unit is
end design_sv_unit;
