library verilog;
use verilog.vl_types.all;
entity lab2_3_tb_sv_unit is
end lab2_3_tb_sv_unit;
