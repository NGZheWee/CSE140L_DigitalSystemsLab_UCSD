library verilog;
use verilog.vl_types.all;
entity lab3_part2_tb is
end lab3_part2_tb;
