library verilog;
use verilog.vl_types.all;
entity light_package is
end light_package;
